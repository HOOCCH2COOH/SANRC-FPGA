// EPCS.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module EPCS (
		input  wire [23:0] addr,          //          addr.addr
		output wire        busy,          //          busy.busy
		input  wire        clkin,         //         clkin.clk
		output wire        data_valid,    //    data_valid.data_valid
		input  wire [7:0]  datain,        //        datain.datain
		output wire [7:0]  dataout,       //       dataout.dataout
		output wire        illegal_write, // illegal_write.illegal_write
		input  wire        rden,          //          rden.rden
		input  wire        read,          //          read.read
		input  wire        reset,         //         reset.reset
		input  wire        wren,          //          wren.wren
		input  wire        write          //         write.write
	);

//	EPCS_asmi_parallel_0 asmi_parallel_0 (
//		.clkin         (clkin),         //         clkin.clk
//		.read          (read),          //          read.read
//		.rden          (rden),          //          rden.rden
//		.addr          (addr),          //          addr.addr
//		.write         (write),         //         write.write
//		.datain        (datain),        //        datain.datain
//		.wren          (wren),          //          wren.wren
//		.reset         (reset),         //         reset.reset
//		.dataout       (dataout),       //       dataout.dataout
//		.busy          (busy),          //          busy.busy
//		.data_valid    (data_valid),    //    data_valid.data_valid
//		.illegal_write (illegal_write)  // illegal_write.illegal_write
//	);

endmodule
